func f(.a(ares), .res(out)); 
endmodule
